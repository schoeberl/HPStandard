-- 
-- Copyright Technical University of Denmark. All rights reserved.
-- This file is part of the Yamp MIPS processor.
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
-- 
--    1. Redistributions of source code must retain the above copyright notice,
--       this list of conditions and the following disclaimer.
-- 
--    2. Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDER ``AS IS'' AND ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES
-- OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN
-- NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF
-- THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation are
-- those of the authors and should not be interpreted as representing official
-- policies, either expressed or implied, of the copyright holder.
-- 


--------------------------------------------------------------------------------
-- Top level of Yamp.
-- Shall be instantiated in an FPGA specific top level.
--
-- Author: Martin Schoeberl (martin@jopdesign.com)
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.yamp_types.all;

entity yamp is
	port(
		clk   : in  std_logic;
		reset : in  std_logic;
		ioout : out io_out_type;
		ioin  : in  io_in_type);
end entity yamp;

architecture rtl of yamp is
	signal feout  : fedec_type;
	signal decout : decex_type;
	signal exout  : exmem_type;
	signal memout : memwb_type;
	signal wbout  : wb_type;

	signal ena : std_logic;

begin
	--	ioout.addr   <= fdout.imm(7 downto 0);
	--	ioout.rd     <= fdout.dec.inp;
	--	ioout.wr     <= fdout.dec.outp;
	--	ioout.wrdata <= exout.accu;

	ena <= '1';                         -- always enabled, no reason to stall (yet)

	fe : entity work.yamp_fetch port map(
			clk, reset, ena, feout
		);
	dec : entity work.yamp_decode port map(
			clk, reset, ena, feout, wbout, decout
		);
	ex : entity work.yamp_execute port map(
			clk, reset, ena, decout, exout
		);
	mem : entity work.yamp_memory port map(
			clk, reset, ena, exout, memout
		);
	wb : entity work.yamp_wback port map(
			clk, reset, ena, memout, wbout
		);

	-- to keep synthesis busy:
	ioout.wrdata <= wbout.rdest.reg.val(15 downto 0);
end;